`timescale 1ns / 1ps

module pe_array(

    );
endmodule
